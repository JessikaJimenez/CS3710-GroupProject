`timescale 1ns/1ns

module tb_datapath #(parameter WIDTH = 16) ();

    reg clk, reset;
    reg pcInstruction, rTypeInstruction;
    reg [1:0] outputSelect;
    reg regWrite, flagSet;
    reg [2:0] aluOp;
    reg pcOverwrite, pcContinue, zeroExtend, luiInstruction;
    wire [WIDTH - 1 : 0] instr; 
    wire [WIDTH - 1 : 0] PC;
    wire [WIDTH - 1 : 0] nextPC;
    wire [WIDTH - 1 : 0] outputFlags;

    datapath #(WIDTH) datpath(
        .clk(clk), 
        .reset(reset), 
        .pcInstruction(pcInstruction), 
        .rTypeInstruction(rTypeInstruction), 
        .outputSelect(outputSelect),
        .regWrite(regWrite), 
        .flagSet(flagSet), 
        .aluOp(aluOp), 
        .pcOverwrite(pcOverwrite), 
        .pcContinue(pcContinue), 
        .zeroExtend(zeroExtend),
        .luiInstruction(luiInstruction), 
        .instr(instr), 
        .PC(PC), 
        .nextPC(nextPC), 
        .outputFlags(outputFlags)
    );
	 
	 
    initial begin
		clk <= 0;
		reset <= 0;
    end
    // Generate clock
    always #10 begin
        clk = ~clk;
    end

endmodule 
