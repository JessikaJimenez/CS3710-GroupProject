// put the address on the LEDs, the read data on one pair of the 7-Segment
// displays, and the write-data on the other pair of 7-segment displays. Use one of
// the pushbuttons to advance the state machine so that we can see each state change.

module memoryFSM ();
  
  
  
  
endmodule
