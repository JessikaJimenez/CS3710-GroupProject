module memoryFSM ();
  
  
  
  
endmodule
