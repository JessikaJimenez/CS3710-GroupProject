// REGISTER FILE MODULE
/*************************************************************/

module RegFile();

endmodule
