// TESTBENCH FOR ALU AND REGISTER FILE
/*************************************************************/

module tb_ALUandRF();

endmodule
