// TOP-LEVEL MODULE
/*************************************************************/

module ALUandRF();

endmodule
